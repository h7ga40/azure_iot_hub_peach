/*
 *		C言語で記述されたアプリケーションから，TECSベースの実行時間分布
 *		集計サービスを呼び出すためのアダプタ用セルタイプの定義
 * 
 *  $Id$
 */
[singleton, active]
celltype tHistogramAdapter {
	call	sHistogram		cHistogram[];
};
