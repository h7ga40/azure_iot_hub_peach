/*
 *		C言語で記述されたアプリケーションから，TECSベースのシステムログ
 *		機能を呼び出すためのアダプタ用セルタイプの定義
 *
 *  $Id$
 */
[singleton, active]
celltype tSysLogAdapter {
	call	sSysLog		cSysLog;
};
